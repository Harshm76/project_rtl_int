packeage top_pkg;
  
  typedef struck {logic [2:0] port_id;
                  logic [11:0] vlan;} connection_addr_t;
  
endpackeage